module sdram_auto_refresh
(
        
);
endmodule